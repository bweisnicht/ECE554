module font_rom_manual(addr,dout);
   input wire [9:0] addr;
   output reg [7:0] dout;
   
   always @(*)
      case(addr)
		   // - 0 - blank
         0:dout = 8'b00000000;
         1:dout = 8'b00000000;
         2:dout = 8'b00000000;
         3:dout = 8'b00000000;
         4:dout = 8'b00000000;
         5:dout = 8'b00000000;
         6:dout = 8'b00000000;
         7:dout = 8'b00000000;
         //" - 1
          8:dout = 8'b11011000;
          9:dout = 8'b11011000;
         10:dout = 8'b11011000;
         11:dout = 8'b00000000;
         12:dout = 8'b00000000;
         13:dout = 8'b00000000;
         14:dout = 8'b00000000;
         15:dout = 8'b00000000;
         //# - 2
         16:dout = 8'b01101100;
         17:dout = 8'b01101100;
         18:dout = 8'b11111110;
         19:dout = 8'b01101100;
         20:dout = 8'b11111110;
         21:dout = 8'b01101100;
         22:dout = 8'b01101100;
         23:dout = 8'b00000000;
         //$ - 3
         24:dout = 8'b00011000;
         25:dout = 8'b01111110;
         26:dout = 8'b11010000;
         27:dout = 8'b01111100;
         28:dout = 8'b00010110;
         29:dout = 8'b11111100;
         30:dout = 8'b00110000;
         31:dout = 8'b00000000;
         //% - 4
         32:dout = 8'b11000000;
         33:dout = 8'b11001100;
         34:dout = 8'b00011000;
         35:dout = 8'b00110000;
         36:dout = 8'b01100000;
         37:dout = 8'b11001100;
         38:dout = 8'b00001100;
         39:dout = 8'b00000000;
         //& - 5
         40:dout = 8'b00011000;
         41:dout = 8'b00110000;
         42:dout = 8'b01100000;
         43:dout = 8'b00000000;
         44:dout = 8'b00000000;
         45:dout = 8'b00000000;
         46:dout = 8'b00000000;
         47:dout = 8'b00000000;
         //` - 6
         48:dout = 8'b00011000;
         49:dout = 8'b00110000;
         50:dout = 8'b01100000;
         51:dout = 8'b00000000;
         52:dout = 8'b00000000;
         53:dout = 8'b00000000;
         54:dout = 8'b00000000;
         55:dout = 8'b00000000;
         //( - 7
         56:dout = 8'b00011000;
         57:dout = 8'b00110000;
         58:dout = 8'b01100000;
         59:dout = 8'b01100000;
         60:dout = 8'b01100000;
         61:dout = 8'b00110000;
         62:dout = 8'b00011000;
         63:dout = 8'b00000000;
         //) - 8
         64:dout = 8'b01100000;
         65:dout = 8'b00110000;
         66:dout = 8'b00011000;
         67:dout = 8'b00011000;
         68:dout = 8'b00011000;
         69:dout = 8'b00110000;
         70:dout = 8'b01100000;
         71:dout = 8'b00000000;
         //* - 9
         72:dout = 8'b00000000;
         73:dout = 8'b00110000;
         74:dout = 8'b11111100;
         75:dout = 8'b01111000;
         76:dout = 8'b11111100;
         77:dout = 8'b00110000;
         78:dout = 8'b00000000;
         79:dout = 8'b00000000;
         //+ - 10
         80:dout = 8'b00000000;
         81:dout = 8'b00110000;
         82:dout = 8'b00110000;
         83:dout = 8'b11111100;
         84:dout = 8'b00110000;
         85:dout = 8'b00110000;
         86:dout = 8'b00000000;
         87:dout = 8'b00000000;
         //; - 11
         88:dout = 8'b00000000;
         89:dout = 8'b00000000;
         90:dout = 8'b00000000;
         91:dout = 8'b00000000;
         92:dout = 8'b00000000;
         93:dout = 8'b00110000;
         94:dout = 8'b00110000;
         95:dout = 8'b01100000;
         //- - 12
         96:dout = 8'b00000000;
         97:dout = 8'b00000000;
         98:dout = 8'b00000000;
         99:dout = 8'b11111100;
         100:dout = 8'b00000000;
         101:dout = 8'b00000000;
         102:dout = 8'b00000000;
         103:dout = 8'b00000000;
         //. - 13
         104:dout = 8'b00000000;
         105:dout = 8'b00000000;
         106:dout = 8'b00000000;
         107:dout = 8'b00000000;
         108:dout = 8'b00000000;
         109:dout = 8'b00110000;
         110:dout = 8'b00110000;
         111:dout = 8'b00000000;
         /// - 14
         112:dout = 8'b00000000;
         113:dout = 8'b00000110;
         114:dout = 8'b00001100;
         115:dout = 8'b00011000;
         116:dout = 8'b00110000;
         117:dout = 8'b01100000;
         118:dout = 8'b11000000;
         119:dout = 8'b00000000;
         //0 - 15
         120:dout = 8'b01111000;
         121:dout = 8'b11001100;
         122:dout = 8'b11011100;
         123:dout = 8'b11111100;
         124:dout = 8'b11101100;
         125:dout = 8'b11001100;
         126:dout = 8'b01111000;
         127:dout = 8'b00000000;
         //1 - 16
         128:dout = 8'b00110000;
         129:dout = 8'b01110000;
         130:dout = 8'b00110000;
         131:dout = 8'b00110000;
         132:dout = 8'b00110000;
         133:dout = 8'b00110000;
         134:dout = 8'b11111100;
         135:dout = 8'b00000000;
         //2 - 17
         136:dout = 8'b01111000;
         137:dout = 8'b11001100;
         138:dout = 8'b00001100;
         139:dout = 8'b00011000;
         140:dout = 8'b00110000;
         141:dout = 8'b01100000;
         142:dout = 8'b11111100;
         143:dout = 8'b00000000;
         //3 - 18
         144:dout = 8'b01111000;
         145:dout = 8'b11001100;
         146:dout = 8'b00001100;
         147:dout = 8'b00111000;
         148:dout = 8'b00001100;
         149:dout = 8'b11001100;
         150:dout = 8'b01111000;
         151:dout = 8'b00000000;
         //4 - 19
         152:dout = 8'b00011000;
         153:dout = 8'b00111000;
         154:dout = 8'b01111000;
         155:dout = 8'b11011000;
         156:dout = 8'b11111100;
         157:dout = 8'b00011000;
         158:dout = 8'b00011000;
         159:dout = 8'b00000000;
         //5 - 20
         160:dout = 8'b11111100;
         161:dout = 8'b11000000;
         162:dout = 8'b11111000;
         163:dout = 8'b00001100;
         164:dout = 8'b00001100;
         165:dout = 8'b11001100;
         166:dout = 8'b01111000;
         167:dout = 8'b00000000;
         //6 - 21
         168:dout = 8'b00111000;
         169:dout = 8'b01100000;
         170:dout = 8'b11000000;
         171:dout = 8'b11111000;
         172:dout = 8'b11001100;
         173:dout = 8'b11001100;
         174:dout = 8'b01111000;
         175:dout = 8'b00000000;
         //7 - 22
         176:dout = 8'b11111100;
         177:dout = 8'b00001100;
         178:dout = 8'b00011000;
         179:dout = 8'b00110000;
         180:dout = 8'b01100000;
         181:dout = 8'b01100000;
         182:dout = 8'b01100000;
         183:dout = 8'b00000000;
         //8 - 23
         184:dout = 8'b01111000;
         185:dout = 8'b11001100;
         186:dout = 8'b11001100;
         187:dout = 8'b01111000;
         188:dout = 8'b11001100;
         189:dout = 8'b11001100;
         190:dout = 8'b01111000;
         191:dout = 8'b00000000;
         //9 - 24
         192:dout = 8'b01111000;
         193:dout = 8'b11001100;
         194:dout = 8'b11001100;
         195:dout = 8'b01111100;
         196:dout = 8'b00001100;
         197:dout = 8'b00011000;
         198:dout = 8'b01110000;
         199:dout = 8'b00000000;
         // - 25
         200:dout = 8'b00000000;
         201:dout = 8'b00000000;
         202:dout = 8'b00110000;
         203:dout = 8'b00110000;
         204:dout = 8'b00000000;
         205:dout = 8'b00110000;
         206:dout = 8'b00110000;
         207:dout = 8'b00000000;
         //// - 26
         208:dout = 8'b00000000;
         209:dout = 8'b00000000;
         210:dout = 8'b00110000;
         211:dout = 8'b00110000;
         212:dout = 8'b00000000;
         213:dout = 8'b00110000;
         214:dout = 8'b00110000;
         215:dout = 8'b01100000;
         //< - 27
         216:dout = 8'b00001100;
         217:dout = 8'b00011000;
         218:dout = 8'b00110000;
         219:dout = 8'b01100000;
         220:dout = 8'b00110000;
         221:dout = 8'b00011000;
         222:dout = 8'b00001100;
         223:dout = 8'b00000000;
         //= - 28
         224:dout = 8'b00000000;
         225:dout = 8'b00000000;
         226:dout = 8'b01111110;
         227:dout = 8'b00000000;
         228:dout = 8'b01111110;
         229:dout = 8'b00000000;
         230:dout = 8'b00000000;
         231:dout = 8'b00000000;
         //> - 29
         232:dout = 8'b01100000;
         233:dout = 8'b00110000;
         234:dout = 8'b00011000;
         235:dout = 8'b00001100;
         236:dout = 8'b00011000;
         237:dout = 8'b00110000;
         238:dout = 8'b01100000;
         239:dout = 8'b00000000;
         //? - 30
         240:dout = 8'b00111100;
         241:dout = 8'b01100110;
         242:dout = 8'b00001100;
         243:dout = 8'b00011000;
         244:dout = 8'b00011000;
         245:dout = 8'b00000000;
         246:dout = 8'b00011000;
         247:dout = 8'b00000000;
         //@ - 31
         248:dout = 8'b01111000;
         249:dout = 8'b11001100;
         250:dout = 8'b11011100;
         251:dout = 8'b11010100;
         252:dout = 8'b11011100;
         253:dout = 8'b11000000;
         254:dout = 8'b01111000;
         255:dout = 8'b00000000;
         //A - 32
         256:dout = 8'b01111000;
         257:dout = 8'b11001100;
         258:dout = 8'b11001100;
         259:dout = 8'b11111100;
         260:dout = 8'b11001100;
         261:dout = 8'b11001100;
         262:dout = 8'b11001100;
         263:dout = 8'b00000000;
         //B - 33
         264:dout = 8'b11111000;
         265:dout = 8'b11001100;
         266:dout = 8'b11001100;
         267:dout = 8'b11111000;
         268:dout = 8'b11001100;
         269:dout = 8'b11001100;
         270:dout = 8'b11111000;
         271:dout = 8'b00000000;
         //C - 34
         272:dout = 8'b01111000;
         273:dout = 8'b11001100;
         274:dout = 8'b11000000;
         275:dout = 8'b11000000;
         276:dout = 8'b11000000;
         277:dout = 8'b11001100;
         278:dout = 8'b01111000;
         279:dout = 8'b00000000;
         //D - 35
         280:dout = 8'b11110000;
         281:dout = 8'b11011000;
         282:dout = 8'b11001100;
         283:dout = 8'b11001100;
         284:dout = 8'b11001100;
         285:dout = 8'b11011000;
         286:dout = 8'b11110000;
         287:dout = 8'b00000000;
         //E - 36
         288:dout = 8'b11111100;
         289:dout = 8'b11000000;
         290:dout = 8'b11000000;
         291:dout = 8'b11111000;
         292:dout = 8'b11000000;
         293:dout = 8'b11000000;
         294:dout = 8'b11111100;
         295:dout = 8'b00000000;
         //F - 37
         296:dout = 8'b11111100;
         297:dout = 8'b11000000;
         298:dout = 8'b11000000;
         299:dout = 8'b11111000;
         300:dout = 8'b11000000;
         301:dout = 8'b11000000;
         302:dout = 8'b11000000;
         303:dout = 8'b00000000;
         //G - 38
         304:dout = 8'b01111000;
         305:dout = 8'b11001100;
         306:dout = 8'b11000000;
         307:dout = 8'b11011100;
         308:dout = 8'b11001100;
         309:dout = 8'b11001100;
         310:dout = 8'b01111000;
         311:dout = 8'b00000000;
         //H - 39
         312:dout = 8'b11001100;
         313:dout = 8'b11001100;
         314:dout = 8'b11001100;
         315:dout = 8'b11111100;
         316:dout = 8'b11001100;
         317:dout = 8'b11001100;
         318:dout = 8'b11001100;
         319:dout = 8'b00000000;
         //I - 40
         320:dout = 8'b11111100;
         321:dout = 8'b00110000;
         322:dout = 8'b00110000;
         323:dout = 8'b00110000;
         324:dout = 8'b00110000;
         325:dout = 8'b00110000;
         326:dout = 8'b11111100;
         327:dout = 8'b00000000;
         //J - 41
         328:dout = 8'b01111100;
         329:dout = 8'b00011000;
         330:dout = 8'b00011000;
         331:dout = 8'b00011000;
         332:dout = 8'b00011000;
         333:dout = 8'b11011000;
         334:dout = 8'b01110000;
         335:dout = 8'b00000000;
         //K - 42
         336:dout = 8'b11001100;
         337:dout = 8'b11011000;
         338:dout = 8'b11110000;
         339:dout = 8'b11100000;
         340:dout = 8'b11110000;
         341:dout = 8'b11011000;
         342:dout = 8'b11001100;
         343:dout = 8'b00000000;
         //L - 43
         344:dout = 8'b11000000;
         345:dout = 8'b11000000;
         346:dout = 8'b11000000;
         347:dout = 8'b11000000;
         348:dout = 8'b11000000;
         349:dout = 8'b11000000;
         350:dout = 8'b11111100;
         351:dout = 8'b00000000;
         //M - 44
         352:dout = 8'b11000110;
         353:dout = 8'b11101110;
         354:dout = 8'b11111110;
         355:dout = 8'b11010110;
         356:dout = 8'b11010110;
         357:dout = 8'b11000110;
         358:dout = 8'b11000110;
         359:dout = 8'b00000000;
         //N - 45
         360:dout = 8'b11001100;
         361:dout = 8'b11001100;
         362:dout = 8'b11101100;
         363:dout = 8'b11111100;
         364:dout = 8'b11011100;
         365:dout = 8'b11001100;
         366:dout = 8'b11001100;
         367:dout = 8'b00000000;
         //O - 46
         368:dout = 8'b01111000;
         369:dout = 8'b11001100;
         370:dout = 8'b11001100;
         371:dout = 8'b11001100;
         372:dout = 8'b11001100;
         373:dout = 8'b11001100;
         374:dout = 8'b01111000;
         375:dout = 8'b00000000;
         //P - 47
         376:dout = 8'b11111000;
         377:dout = 8'b11001100;
         378:dout = 8'b11001100;
         379:dout = 8'b11111000;
         380:dout = 8'b11000000;
         381:dout = 8'b11000000;
         382:dout = 8'b11000000;
         383:dout = 8'b00000000;
         //Q - 48
         384:dout = 8'b01111000;
         385:dout = 8'b11001100;
         386:dout = 8'b11001100;
         387:dout = 8'b11001100;
         388:dout = 8'b11010100;
         389:dout = 8'b11011000;
         390:dout = 8'b01101100;
         391:dout = 8'b00000000;
         //R - 49
         392:dout = 8'b11111000;
         393:dout = 8'b11001100;
         394:dout = 8'b11001100;
         395:dout = 8'b11111000;
         396:dout = 8'b11011000;
         397:dout = 8'b11001100;
         398:dout = 8'b11001100;
         399:dout = 8'b00000000;
         //S - 50
         400:dout = 8'b01111000;
         401:dout = 8'b11001100;
         402:dout = 8'b11000000;
         403:dout = 8'b01111100;
         404:dout = 8'b00001100;
         405:dout = 8'b11001100;
         406:dout = 8'b01111000;
         407:dout = 8'b00000000;
         //T - 51
         408:dout = 8'b11111100;
         409:dout = 8'b00110000;
         410:dout = 8'b00110000;
         411:dout = 8'b00110000;
         412:dout = 8'b00110000;
         413:dout = 8'b00110000;
         414:dout = 8'b00110000;
         415:dout = 8'b00000000;
         //U - 52
         416:dout = 8'b11001100;
         417:dout = 8'b11001100;
         418:dout = 8'b11001100;
         419:dout = 8'b11001100;
         420:dout = 8'b11001100;
         421:dout = 8'b11001100;
         422:dout = 8'b01111000;
         423:dout = 8'b00000000;
         //V - 53
         424:dout = 8'b11001100;
         425:dout = 8'b11001100;
         426:dout = 8'b11001100;
         427:dout = 8'b11001100;
         428:dout = 8'b11001100;
         429:dout = 8'b01111000;
         430:dout = 8'b00110000;
         431:dout = 8'b00000000;
         //W - 54
         432:dout = 8'b11000110;
         433:dout = 8'b11000110;
         434:dout = 8'b11010110;
         435:dout = 8'b11010110;
         436:dout = 8'b11111110;
         437:dout = 8'b11101110;
         438:dout = 8'b11001100;
         439:dout = 8'b00000000;
         //X - 55
         440:dout = 8'b11001100;
         441:dout = 8'b11001100;
         442:dout = 8'b01111000;
         443:dout = 8'b00110000;
         444:dout = 8'b01111000;
         445:dout = 8'b11001100;
         446:dout = 8'b11001100;
         447:dout = 8'b00000000;
         //Y - 56
         448:dout = 8'b11001100;
         449:dout = 8'b11001100;
         450:dout = 8'b11001100;
         451:dout = 8'b01111000;
         452:dout = 8'b00110000;
         453:dout = 8'b00110000;
         454:dout = 8'b00110000;
         455:dout = 8'b00000000;
         //Z - 57
         456:dout = 8'b11111100;
         457:dout = 8'b00001100;
         458:dout = 8'b00011000;
         459:dout = 8'b00110000;
         460:dout = 8'b01100000;
         461:dout = 8'b11000000;
         462:dout = 8'b11111100;
         463:dout = 8'b00000000;
         //[ - 58
         464:dout = 8'b11111000;
         465:dout = 8'b11000000;
         466:dout = 8'b11000000;
         467:dout = 8'b11000000;
         468:dout = 8'b11000000;
         469:dout = 8'b11000000;
         470:dout = 8'b11111000;
         471:dout = 8'b00000000;
         //\ - 59
         472:dout = 8'b00000000;
         473:dout = 8'b01100000;
         474:dout = 8'b00110000;
         475:dout = 8'b00011000;
         476:dout = 8'b00001100;
         477:dout = 8'b00000110;
         478:dout = 8'b00000000;
         479:dout = 8'b00000000;
         //] - 60
         480:dout = 8'b01111100;
         481:dout = 8'b00001100;
         482:dout = 8'b00001100;
         483:dout = 8'b00001100;
         484:dout = 8'b00001100;
         485:dout = 8'b00001100;
         486:dout = 8'b01111100;
         487:dout = 8'b00000000;
         //^ - 61
         488:dout = 8'b00110000;
         489:dout = 8'b01111000;
         490:dout = 8'b11001100;
         491:dout = 8'b10000100;
         492:dout = 8'b00000000;
         493:dout = 8'b00000000;
         494:dout = 8'b00000000;
         495:dout = 8'b00000000;
         //_ - 62
         496:dout = 8'b00000000;
         497:dout = 8'b00000000;
         498:dout = 8'b00000000;
         499:dout = 8'b00000000;
         500:dout = 8'b00000000;
         501:dout = 8'b00000000;
         502:dout = 8'b00000000;
         503:dout = 8'b11111111;
         //GBP - 63
         504:dout = 8'b00110000;
         505:dout = 8'b01101100;
         506:dout = 8'b01100000;
         507:dout = 8'b11111000;
         508:dout = 8'b01100000;
         509:dout = 8'b01100000;
         510:dout = 8'b11111100;
         511:dout = 8'b00000000;
         //a - 64
         512:dout = 8'b00000000;
         513:dout = 8'b00000000;
         514:dout = 8'b01111000;
         515:dout = 8'b00001100;
         516:dout = 8'b01111100;
         517:dout = 8'b11001100;
         518:dout = 8'b01111100;
         519:dout = 8'b00000000;
         //b - 65
         520:dout = 8'b11000000;
         521:dout = 8'b11000000;
         522:dout = 8'b11111000;
         523:dout = 8'b11001100;
         524:dout = 8'b11001100;
         525:dout = 8'b11001100;
         526:dout = 8'b11111000;
         527:dout = 8'b00000000;
         //c - 66
         528:dout = 8'b00000000;
         529:dout = 8'b00000000;
         530:dout = 8'b01111000;
         531:dout = 8'b11001100;
         532:dout = 8'b11000000;
         533:dout = 8'b11001100;
         534:dout = 8'b01111000;
         535:dout = 8'b00000000;
         //d - 67
         536:dout = 8'b00001100;
         537:dout = 8'b00001100;
         538:dout = 8'b01111100;
         539:dout = 8'b11001100;
         540:dout = 8'b11001100;
         541:dout = 8'b11001100;
         542:dout = 8'b01111100;
         543:dout = 8'b00000000;
         //e - 68
         544:dout = 8'b00000000;
         545:dout = 8'b00000000;
         546:dout = 8'b01111000;
         547:dout = 8'b11001100;
         548:dout = 8'b11111100;
         549:dout = 8'b11000000;
         550:dout = 8'b01111000;
         551:dout = 8'b00000000;
         //f - 69
         552:dout = 8'b00111000;
         553:dout = 8'b01100000;
         554:dout = 8'b01100000;
         555:dout = 8'b11111000;
         556:dout = 8'b01100000;
         557:dout = 8'b01100000;
         558:dout = 8'b01100000;
         559:dout = 8'b00000000;
         //g - 70
         560:dout = 8'b00000000;
         561:dout = 8'b00000000;
         562:dout = 8'b01111100;
         563:dout = 8'b11001100;
         564:dout = 8'b11001100;
         565:dout = 8'b01111100;
         566:dout = 8'b00001100;
         567:dout = 8'b00111000;
         //h - 71
         568:dout = 8'b11000000;
         569:dout = 8'b11000000;
         570:dout = 8'b11111000;
         571:dout = 8'b11001100;
         572:dout = 8'b11001100;
         573:dout = 8'b11001100;
         574:dout = 8'b11001100;
         575:dout = 8'b00000000;
         //i - 72
         576:dout = 8'b00110000;
         577:dout = 8'b00000000;
         578:dout = 8'b01110000;
         579:dout = 8'b00110000;
         580:dout = 8'b00110000;
         581:dout = 8'b00110000;
         582:dout = 8'b01111000;
         583:dout = 8'b00000000;
         //j - 73
         584:dout = 8'b00110000;
         585:dout = 8'b00000000;
         586:dout = 8'b01110000;
         587:dout = 8'b00110000;
         588:dout = 8'b00110000;
         589:dout = 8'b00110000;
         590:dout = 8'b00110000;
         591:dout = 8'b11100000;
         //k - 74
         592:dout = 8'b11000000;
         593:dout = 8'b11000000;
         594:dout = 8'b11001100;
         595:dout = 8'b11011000;
         596:dout = 8'b11110000;
         597:dout = 8'b11011000;
         598:dout = 8'b11001100;
         599:dout = 8'b00000000;
         //l - 75
         600:dout = 8'b11100000;
         601:dout = 8'b01100000;
         602:dout = 8'b01100000;
         603:dout = 8'b01100000;
         604:dout = 8'b01100000;
         605:dout = 8'b01100000;
         606:dout = 8'b11110000;
         607:dout = 8'b00000000;
         //m - 76
         608:dout = 8'b00000000;
         609:dout = 8'b00000000;
         610:dout = 8'b01101100;
         611:dout = 8'b11111110;
         612:dout = 8'b11010110;
         613:dout = 8'b11010110;
         614:dout = 8'b11000110;
         615:dout = 8'b00000000;
         //n - 77
         616:dout = 8'b00000000;
         617:dout = 8'b00000000;
         618:dout = 8'b11111000;
         619:dout = 8'b11001100;
         620:dout = 8'b11001100;
         621:dout = 8'b11001100;
         622:dout = 8'b11001100;
         623:dout = 8'b00000000;
         //o - 78
         624:dout = 8'b00000000;
         625:dout = 8'b00000000;
         626:dout = 8'b01111000;
         627:dout = 8'b11001100;
         628:dout = 8'b11001100;
         629:dout = 8'b11001100;
         630:dout = 8'b01111000;
         631:dout = 8'b00000000;
         //p - 79
         632:dout = 8'b00000000;
         633:dout = 8'b00000000;
         634:dout = 8'b11111000;
         635:dout = 8'b11001100;
         636:dout = 8'b11001100;
         637:dout = 8'b11111000;
         638:dout = 8'b11000000;
         639:dout = 8'b11000000;
         //q - 80
         640:dout = 8'b00000000;
         641:dout = 8'b00000000;
         642:dout = 8'b01111100;
         643:dout = 8'b11001100;
         644:dout = 8'b11001100;
         645:dout = 8'b01111100;
         646:dout = 8'b00001100;
         647:dout = 8'b00001110;
         //r - 81
         648:dout = 8'b00000000;
         649:dout = 8'b00000000;
         650:dout = 8'b11011000;
         651:dout = 8'b11101100;
         652:dout = 8'b11000000;
         653:dout = 8'b11000000;
         654:dout = 8'b11000000;
         655:dout = 8'b00000000;
         //s - 82
         656:dout = 8'b00000000;
         657:dout = 8'b00000000;
         658:dout = 8'b01111100;
         659:dout = 8'b11000000;
         660:dout = 8'b01111000;
         661:dout = 8'b00001100;
         662:dout = 8'b11111000;
         663:dout = 8'b00000000;
         //t - 83
         664:dout = 8'b01100000;
         665:dout = 8'b01100000;
         666:dout = 8'b11111000;
         667:dout = 8'b01100000;
         668:dout = 8'b01100000;
         669:dout = 8'b01100000;
         670:dout = 8'b00111000;
         671:dout = 8'b00000000;
         //u - 84
         672:dout = 8'b00000000;
         673:dout = 8'b00000000;
         674:dout = 8'b11001100;
         675:dout = 8'b11001100;
         676:dout = 8'b11001100;
         677:dout = 8'b11001100;
         678:dout = 8'b01111100;
         679:dout = 8'b00000000;
         //v - 85
         680:dout = 8'b00000000;
         681:dout = 8'b00000000;
         682:dout = 8'b11001100;
         683:dout = 8'b11001100;
         684:dout = 8'b11001100;
         685:dout = 8'b01111000;
         686:dout = 8'b00110000;
         687:dout = 8'b00000000;
         //w - 86
         688:dout = 8'b00000000;
         689:dout = 8'b00000000;
         690:dout = 8'b11000110;
         691:dout = 8'b11010110;
         692:dout = 8'b11010110;
         693:dout = 8'b11111110;
         694:dout = 8'b01101100;
         695:dout = 8'b00000000;
         //x - 87
         696:dout = 8'b00000000;
         697:dout = 8'b00000000;
         698:dout = 8'b11001100;
         699:dout = 8'b01111000;
         700:dout = 8'b00110000;
         701:dout = 8'b01111000;
         702:dout = 8'b11001100;
         703:dout = 8'b00000000;
         //y - 88
         704:dout = 8'b00000000;
         705:dout = 8'b00000000;
         706:dout = 8'b11001100;
         707:dout = 8'b11001100;
         708:dout = 8'b11001100;
         709:dout = 8'b01111100;
         710:dout = 8'b00001100;
         711:dout = 8'b01111000;
         //z - 89
         712:dout = 8'b00000000;
         713:dout = 8'b00000000;
         714:dout = 8'b11111100;
         715:dout = 8'b00011000;
         716:dout = 8'b00110000;
         717:dout = 8'b01100000;
         718:dout = 8'b11111100;
         719:dout = 8'b00000000;
         //{ - 90
         720:dout = 8'b00001100;
         721:dout = 8'b00011000;
         722:dout = 8'b00011000;
         723:dout = 8'b01110000;
         724:dout = 8'b00011000;
         725:dout = 8'b00011000;
         726:dout = 8'b00001100;
         727:dout = 8'b00000000;
         //| - 91
         728:dout = 8'b00011000;
         729:dout = 8'b00011000;
         730:dout = 8'b00011000;
         731:dout = 8'b00000000;
         732:dout = 8'b00011000;
         733:dout = 8'b00011000;
         734:dout = 8'b00011000;
         735:dout = 8'b00000000;
         //} - 92
         736:dout = 8'b01100000;
         737:dout = 8'b00110000;
         738:dout = 8'b00110000;
         739:dout = 8'b00011100;
         740:dout = 8'b00110000;
         741:dout = 8'b00110000;
         742:dout = 8'b01100000;
         743:dout = 8'b00000000;
		   // ! - 93
         744:dout = 8'b00110000;
         745:dout = 8'b00110000;
         746:dout = 8'b00110000;
         747:dout = 8'b00110000;
         748:dout = 8'b00110000;
         749:dout = 8'b00000000;
         750:dout = 8'b00110000;
         751:dout = 8'b00000000;
         // - 94 - left blank
         752:dout = 8'b00000000;
         753:dout = 8'b00000000;
         754:dout = 8'b00000000;
         755:dout = 8'b00000000;
         756:dout = 8'b00000000;
         757:dout = 8'b00000000;
         758:dout = 8'b00000000;
         759:dout = 8'b00000000;
         // - 95 - left blank
         760:dout = 8'b00000000;
         761:dout = 8'b00000000;
         762:dout = 8'b00000000;
         763:dout = 8'b00000000;
         764:dout = 8'b00000000;
         765:dout = 8'b00000000;
         766:dout = 8'b00000000;
         767:dout = 8'b00000000;
         // - 96 - Column cap beginning
         768:dout = 8'b10000000;
         769:dout = 8'b10000000;
         770:dout = 8'b10000000;
         771:dout = 8'b10000000;
         772:dout = 8'b10000000;
         773:dout = 8'b10000000;
         774:dout = 8'b10000000;
         775:dout = 8'b10000000;
         // - 97
         776:dout = 8'b11000000;
         777:dout = 8'b11000000;
         778:dout = 8'b11000000;
         779:dout = 8'b11000000;
         780:dout = 8'b11000000;
         781:dout = 8'b11000000;
         782:dout = 8'b11000000;
         783:dout = 8'b11000000;
         // - 98
         784:dout = 8'b11100000;
         785:dout = 8'b11100000;
         786:dout = 8'b11100000;
         787:dout = 8'b11100000;
         788:dout = 8'b11100000;
         789:dout = 8'b11100000;
         790:dout = 8'b11100000;
         791:dout = 8'b11100000;
         // - 99
         792:dout = 8'b11110000;
         793:dout = 8'b11110000;
         794:dout = 8'b11110000;
         795:dout = 8'b11110000;
         796:dout = 8'b11110000;
         797:dout = 8'b11110000;
         798:dout = 8'b11110000;
         799:dout = 8'b11110000;
         // - 100
         800:dout = 8'b11111000;
         801:dout = 8'b11111000;
         802:dout = 8'b11111000;
         803:dout = 8'b11111000;
         804:dout = 8'b11111000;
         805:dout = 8'b11111000;
         806:dout = 8'b11111000;
         807:dout = 8'b11111000;
         // - 101
         808:dout = 8'b11111100;
         809:dout = 8'b11111100;
         810:dout = 8'b11111100;
         811:dout = 8'b11111100;
         812:dout = 8'b11111100;
         813:dout = 8'b11111100;
         814:dout = 8'b11111100;
         815:dout = 8'b11111100;
         // - 102
         816:dout = 8'b11111110;
         817:dout = 8'b11111110;
         818:dout = 8'b11111110;
         819:dout = 8'b11111110;
         820:dout = 8'b11111110;
         821:dout = 8'b11111110;
         822:dout = 8'b11111110;
         823:dout = 8'b11111110;
         // - 103 - Column block
         824:dout = 8'b11111111;
         825:dout = 8'b11111111;
         826:dout = 8'b11111111;
         827:dout = 8'b11111111;
         828:dout = 8'b11111111;
         829:dout = 8'b11111111;
         830:dout = 8'b11111111;
         831:dout = 8'b11111111;
         // - 104
         832:dout = 8'b01111111;
         833:dout = 8'b01111111;
         834:dout = 8'b01111111;
         835:dout = 8'b01111111;
         836:dout = 8'b01111111;
         837:dout = 8'b01111111;
         838:dout = 8'b01111111;
         839:dout = 8'b01111111;
         // - 105
         840:dout = 8'b00111111;
         841:dout = 8'b00111111;
         842:dout = 8'b00111111;
         843:dout = 8'b00111111;
         844:dout = 8'b00111111;
         845:dout = 8'b00111111;
         846:dout = 8'b00111111;
         847:dout = 8'b00111111;
         // - 106
         848:dout = 8'b00011111;
         849:dout = 8'b00011111;
         850:dout = 8'b00011111;
         851:dout = 8'b00011111;
         852:dout = 8'b00011111;
         853:dout = 8'b00011111;
         854:dout = 8'b00011111;
         855:dout = 8'b00011111;
         // - 107
         856:dout = 8'b00001111;
         857:dout = 8'b00001111;
         858:dout = 8'b00001111;
         859:dout = 8'b00001111;
         860:dout = 8'b00001111;
         861:dout = 8'b00001111;
         862:dout = 8'b00001111;
         863:dout = 8'b00001111;
         // - 108
         864:dout = 8'b00000111;
         865:dout = 8'b00000111;
         866:dout = 8'b00000111;
         867:dout = 8'b00000111;
         868:dout = 8'b00000111;
         869:dout = 8'b00000111;
         870:dout = 8'b00000111;
         871:dout = 8'b00000111;
         // - 109
         872:dout = 8'b00000011;
         873:dout = 8'b00000011;
         874:dout = 8'b00000011;
         875:dout = 8'b00000011;
         876:dout = 8'b00000011;
         877:dout = 8'b00000011;
         878:dout = 8'b00000011;
         879:dout = 8'b00000011;
         // - 110 - Column base ending
         880:dout = 8'b00000001; 
         881:dout = 8'b00000001;
         882:dout = 8'b00000001;
         883:dout = 8'b00000001;
         884:dout = 8'b00000001;
         885:dout = 8'b00000001;
         886:dout = 8'b00000001;
         887:dout = 8'b00000001;
         // - 111
         888:dout = 8'b00011000;
         889:dout = 8'b00011000;
         890:dout = 8'b00011000;
         891:dout = 8'b00011000;
         892:dout = 8'b00011000;
         893:dout = 8'b00011000;
         894:dout = 8'b00011000;
         895:dout = 8'b00011000;
         // - 112
         896:dout = 8'b00000000;
         897:dout = 8'b00000000;
         898:dout = 8'b00000000;
         899:dout = 8'b11111111; 
         900:dout = 8'b11111111; 
         901:dout = 8'b00000000;
         902:dout = 8'b00000000;
         903:dout = 8'b00000000;
         // - 113
         904:dout = 8'b00011000;
         905:dout = 8'b00011000;
         906:dout = 8'b00011000;
         907:dout = 8'b11111111; 
         908:dout = 8'b11111111; 
         909:dout = 8'b00011000;
         910:dout = 8'b00011000;
         911:dout = 8'b00011000;
         // - 114
         912:dout = 8'b00011000;
         913:dout = 8'b00011000;
         914:dout = 8'b00011000;
         915:dout = 8'b11111000; 
         916:dout = 8'b11111000; 
         917:dout = 8'b00000000;
         918:dout = 8'b00000000;
         919:dout = 8'b00000000;
         // - 115
         920:dout = 8'b00011000;
         921:dout = 8'b00011000;
         922:dout = 8'b00011000;
         923:dout = 8'b00011111; 
         924:dout = 8'b00011111; 
         925:dout = 8'b00000000;
         926:dout = 8'b00000000;
         927:dout = 8'b00000000;
         // - 116
         928:dout = 8'b00000000;
         929:dout = 8'b00000000;
         930:dout = 8'b00000000;
         931:dout = 8'b11111000; 
         932:dout = 8'b11111000; 
         933:dout = 8'b00011000;
         934:dout = 8'b00011000;
         935:dout = 8'b00011000;
         // - 117
         936:dout = 8'b00000000;
         937:dout = 8'b00000000;
         938:dout = 8'b00000000;
         939:dout = 8'b00011111; 
         940:dout = 8'b00011111; 
         941:dout = 8'b00011000;
         942:dout = 8'b00011000;
         943:dout = 8'b00011000;
         // - 118
         944:dout = 8'b00011000;
         945:dout = 8'b00011000;
         946:dout = 8'b00011000;
         947:dout = 8'b11111000; 
         948:dout = 8'b11111000; 
         949:dout = 8'b00011000;
         950:dout = 8'b00011000;
         951:dout = 8'b00011000;
         // - 119
         952:dout = 8'b00011000;
         953:dout = 8'b00011000;
         954:dout = 8'b00011000;
         955:dout = 8'b00011111; 
         956:dout = 8'b00011111; 
         957:dout = 8'b00011000;
         958:dout = 8'b00011000;
         959:dout = 8'b00011000;
         // - 120
         960:dout = 8'b00000000;
         961:dout = 8'b00000000;
         962:dout = 8'b00000000;
         963:dout = 8'b11111111; 
         964:dout = 8'b11111111; 
         965:dout = 8'b00011000;
         966:dout = 8'b00011000;
         967:dout = 8'b00011000;
         // - 121
         968:dout = 8'b00011000;
         969:dout = 8'b00011000;
         970:dout = 8'b00011000;
         971:dout = 8'b11111111; 
         972:dout = 8'b11111111; 
         973:dout = 8'b00000000;
         974:dout = 8'b00000000;
         975:dout = 8'b00000000;
         // - 122
         976:dout = 8'b00000000;
         977:dout = 8'b00000000;
         978:dout = 8'b00000000;
         979:dout = 8'b00011000;
         980:dout = 8'b00011000;
         981:dout = 8'b00000000;
         982:dout = 8'b00000000;
         983:dout = 8'b00000000;
         //... - 123
         984:dout = 8'b00000000;
         985:dout = 8'b00000000;
         986:dout = 8'b00000000;
         987:dout = 8'b00000000;
         988:dout = 8'b00000000;
         989:dout = 8'b01010100;
         990:dout = 8'b01010100;
         991:dout = 8'b00000000;
         // - 124
         992:dout = 8'b01010101;
         993:dout = 8'b10101010;
         994:dout = 8'b01010101;
         995:dout = 8'b10101010;
         996:dout = 8'b01010101;
         997:dout = 8'b10101010;
         998:dout = 8'b01010101;
         999:dout = 8'b10101010;
         // - 125
         1000:dout = 8'b10101010;
         1001:dout = 8'b01010101;
         1002:dout = 8'b10101010;
         1003:dout = 8'b01010101;
         1004:dout = 8'b10101010;
         1005:dout = 8'b01010101;
         1006:dout = 8'b10101010;
         1007:dout = 8'b01010101;
         // - 126
         1008:dout = 8'b10101010;
         1009:dout = 8'b10101010;
         1010:dout = 8'b10101010;
         1011:dout = 8'b10101010;
         1012:dout = 8'b10101010;
         1013:dout = 8'b10101010;
         1014:dout = 8'b10101010;
         1015:dout = 8'b10101010;
         // - 127
         1016:dout = 8'b01010101;
         1017:dout = 8'b01010101;
         1018:dout = 8'b01010101;
         1019:dout = 8'b01010101;
         1020:dout = 8'b01010101;
         1021:dout = 8'b01010101;
         1022:dout = 8'b01010101;
         1023:dout = 8'b01010101;
      endcase
endmodule
